`timescale 1ns / 1ps

module BROM(
	input	[7:1]	adr_i,
	input		stb_i,
	output		ack_o,
	output	[15:0]	dat_o
);
	reg	[15:0]	dat_o;
	assign ack_o = stb_i;
	always @(*) begin
		case(adr_i)
		7'd0: dat_o = 16'h0113;
		7'd1: dat_o = 16'h0000;
		7'd2: dat_o = 16'h01B7;
		7'd3: dat_o = 16'h0010;
		7'd4: dat_o = 16'h0113;
		7'd5: dat_o = 16'h0011;
		7'd6: dat_o = 16'h5213;
		7'd7: dat_o = 16'h0101;
		7'd8: dat_o = 16'h9123;
		7'd9: dat_o = 16'h0041;
		7'd10: dat_o = 16'hF06F;
		7'd11: dat_o = 16'hFF5F;
		7'd12: dat_o = 16'hCCCC;
		7'd13: dat_o = 16'hCCCC;
		7'd14: dat_o = 16'hCCCC;
		7'd15: dat_o = 16'hCCCC;
		7'd16: dat_o = 16'hCCCC;
		7'd17: dat_o = 16'hCCCC;
		7'd18: dat_o = 16'hCCCC;
		7'd19: dat_o = 16'hCCCC;
		7'd20: dat_o = 16'hCCCC;
		7'd21: dat_o = 16'hCCCC;
		7'd22: dat_o = 16'hCCCC;
		7'd23: dat_o = 16'hCCCC;
		7'd24: dat_o = 16'hCCCC;
		7'd25: dat_o = 16'hCCCC;
		7'd26: dat_o = 16'hCCCC;
		7'd27: dat_o = 16'hCCCC;
		7'd28: dat_o = 16'hCCCC;
		7'd29: dat_o = 16'hCCCC;
		7'd30: dat_o = 16'hCCCC;
		7'd31: dat_o = 16'hCCCC;
		7'd32: dat_o = 16'hCCCC;
		7'd33: dat_o = 16'hCCCC;
		7'd34: dat_o = 16'hCCCC;
		7'd35: dat_o = 16'hCCCC;
		7'd36: dat_o = 16'hCCCC;
		7'd37: dat_o = 16'hCCCC;
		7'd38: dat_o = 16'hCCCC;
		7'd39: dat_o = 16'hCCCC;
		7'd40: dat_o = 16'hCCCC;
		7'd41: dat_o = 16'hCCCC;
		7'd42: dat_o = 16'hCCCC;
		7'd43: dat_o = 16'hCCCC;
		7'd44: dat_o = 16'hCCCC;
		7'd45: dat_o = 16'hCCCC;
		7'd46: dat_o = 16'hCCCC;
		7'd47: dat_o = 16'hCCCC;
		7'd48: dat_o = 16'hCCCC;
		7'd49: dat_o = 16'hCCCC;
		7'd50: dat_o = 16'hCCCC;
		7'd51: dat_o = 16'hCCCC;
		7'd52: dat_o = 16'hCCCC;
		7'd53: dat_o = 16'hCCCC;
		7'd54: dat_o = 16'hCCCC;
		7'd55: dat_o = 16'hCCCC;
		7'd56: dat_o = 16'hCCCC;
		7'd57: dat_o = 16'hCCCC;
		7'd58: dat_o = 16'hCCCC;
		7'd59: dat_o = 16'hCCCC;
		7'd60: dat_o = 16'hCCCC;
		7'd61: dat_o = 16'hCCCC;
		7'd62: dat_o = 16'hCCCC;
		7'd63: dat_o = 16'hCCCC;
		7'd64: dat_o = 16'hCCCC;
		7'd65: dat_o = 16'hCCCC;
		7'd66: dat_o = 16'hCCCC;
		7'd67: dat_o = 16'hCCCC;
		7'd68: dat_o = 16'hCCCC;
		7'd69: dat_o = 16'hCCCC;
		7'd70: dat_o = 16'hCCCC;
		7'd71: dat_o = 16'hCCCC;
		7'd72: dat_o = 16'hCCCC;
		7'd73: dat_o = 16'hCCCC;
		7'd74: dat_o = 16'hCCCC;
		7'd75: dat_o = 16'hCCCC;
		7'd76: dat_o = 16'hCCCC;
		7'd77: dat_o = 16'hCCCC;
		7'd78: dat_o = 16'hCCCC;
		7'd79: dat_o = 16'hCCCC;
		7'd80: dat_o = 16'hCCCC;
		7'd81: dat_o = 16'hCCCC;
		7'd82: dat_o = 16'hCCCC;
		7'd83: dat_o = 16'hCCCC;
		7'd84: dat_o = 16'hCCCC;
		7'd85: dat_o = 16'hCCCC;
		7'd86: dat_o = 16'hCCCC;
		7'd87: dat_o = 16'hCCCC;
		7'd88: dat_o = 16'hCCCC;
		7'd89: dat_o = 16'hCCCC;
		7'd90: dat_o = 16'hCCCC;
		7'd91: dat_o = 16'hCCCC;
		7'd92: dat_o = 16'hCCCC;
		7'd93: dat_o = 16'hCCCC;
		7'd94: dat_o = 16'hCCCC;
		7'd95: dat_o = 16'hCCCC;
		7'd96: dat_o = 16'hCCCC;
		7'd97: dat_o = 16'hCCCC;
		7'd98: dat_o = 16'hCCCC;
		7'd99: dat_o = 16'hCCCC;
		7'd100: dat_o = 16'hCCCC;
		7'd101: dat_o = 16'hCCCC;
		7'd102: dat_o = 16'hCCCC;
		7'd103: dat_o = 16'hCCCC;
		7'd104: dat_o = 16'hCCCC;
		7'd105: dat_o = 16'hCCCC;
		7'd106: dat_o = 16'hCCCC;
		7'd107: dat_o = 16'hCCCC;
		7'd108: dat_o = 16'hCCCC;
		7'd109: dat_o = 16'hCCCC;
		7'd110: dat_o = 16'hCCCC;
		7'd111: dat_o = 16'hCCCC;
		7'd112: dat_o = 16'hCCCC;
		7'd113: dat_o = 16'hCCCC;
		7'd114: dat_o = 16'hCCCC;
		7'd115: dat_o = 16'hCCCC;
		7'd116: dat_o = 16'hCCCC;
		7'd117: dat_o = 16'hCCCC;
		7'd118: dat_o = 16'hCCCC;
		7'd119: dat_o = 16'hCCCC;
		7'd120: dat_o = 16'hCCCC;
		7'd121: dat_o = 16'hCCCC;
		7'd122: dat_o = 16'hCCCC;
		7'd123: dat_o = 16'hCCCC;
		7'd124: dat_o = 16'hCCCC;
		7'd125: dat_o = 16'hCCCC;
		7'd126: dat_o = 16'hCCCC;
		7'd127: dat_o = 16'hCCCC;
		endcase
	end
endmodule
